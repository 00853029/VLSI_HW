module top(
    input  logic           cpu_clk,
    input  logic           axi_clk,
    input  logic           rom_clk,
    input  logic           dram_clk,
    input  logic           sram_clk,
    input  logic           cpu_rst,
    input  logic           axi_rst,
    input  logic           rom_rst,
    input  logic           dram_rst,
    input  logic           sram_rst,
    input  logic           sensor_ready,
    input  logic [   31:0] sensor_out,
    output logic           sensor_en,
    input  logic [   31:0] ROM_out,
    input  logic [   31:0] DRAM_Q,
    output logic           ROM_read,
    output logic           ROM_enable,
    output logic [   11:0] ROM_address,
    output logic           DRAM_CSn,
    output logic [    3:0] DRAM_WEn,
    output logic           DRAM_RASn,
    output logic           DRAM_CASn,
    output logic [   10:0] DRAM_A,
    output logic [   31:0] DRAM_D,
    input  logic           DRAM_valid
);



endmodule


